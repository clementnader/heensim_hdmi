----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/05/2021 12:07:46 PM
-- Package Name: neurons_platform_spec_pkg
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;


package neurons_platform_spec_pkg is
    
    constant C_PLATFORM_NAME : STRING := "ZedBoard";
    
end package;


package body neurons_platform_spec_pkg is
    
end package body;
